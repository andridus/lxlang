module compiler

enum Identifier {
	x
	y
	atom
	integer
	nil
	f
	string
	extfunc
	list
	commands
	float
	fr
	field_flags
	alloc
	literal
}
