module compiler

fn test_extract_vars() {
	assert true
}
