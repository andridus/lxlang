module erl

const max_u8 = 255
const max_u16 = 65535
const max_u32 = u64(4294967295)
const max_u64 = u64(18446744073709551615)
const max_i8 = 127
const max_i6 = 32767
const max_i32 = u64(2147483647)
const max_i64 = u64(9223372036854775807)
